MACRO block_126x981_68
   SIZE 47.88 BY 186.39 ;
END block_126x981_68

MACRO block_533x4743_849
   SIZE 202.54 BY 901.17 ;
END block_533x4743_849

MACRO block_416x441_106
   SIZE 158.08 BY 83.79 ;
END block_416x441_106

MACRO block_1024x1296_101
   SIZE 389.12 BY 246.24 ;
END block_1024x1296_101

MACRO block_341x369_78
   SIZE 129.58 BY 70.11 ;
END block_341x369_78

MACRO block_533x1791_321
   SIZE 202.54 BY 340.29 ;
END block_533x1791_321

MACRO block_779x3546_628
   SIZE 296.02 BY 673.74 ;
END block_779x3546_628

MACRO block_416x441_108
   SIZE 158.08 BY 83.79 ;
END block_416x441_108

MACRO block_1829x2628_275
   SIZE 695.02 BY 499.32 ;
END block_1829x2628_275

MACRO block_341x369_84
   SIZE 129.58 BY 70.11 ;
END block_341x369_84

MACRO block_1338x2115_224
   SIZE 508.44 BY 401.85 ;
END block_1338x2115_224

MACRO block_341x369_82
   SIZE 129.58 BY 70.11 ;
END block_341x369_82

MACRO block_1338x2799_288
   SIZE 508.44 BY 531.81 ;
END block_1338x2799_288

MACRO block_546x675_103
   SIZE 207.48 BY 128.25 ;
END block_546x675_103

MACRO block_4656x6120_609
   SIZE 1769.28 BY 1162.8 ;
END block_4656x6120_609

MACRO block_646x2655_74
   SIZE 245.48 BY 504.45 ;
END block_646x2655_74

MACRO block_779x2529_460
   SIZE 296.02 BY 480.51 ;
END block_779x2529_460

MACRO block_341x369_80
   SIZE 129.58 BY 70.11 ;
END block_341x369_80

MACRO block_1338x4491_807
   SIZE 508.44 BY 853.29 ;
END block_1338x4491_807

MACRO block_416x441_110
   SIZE 158.08 BY 83.79 ;
END block_416x441_110

MACRO block_1338x6147_608
   SIZE 508.44 BY 1167.93 ;
END block_1338x6147_608

MACRO block_416x441_118
   SIZE 158.08 BY 83.79 ;
END block_416x441_118

MACRO block_779x1467_106
   SIZE 296.02 BY 278.73 ;
END block_779x1467_106

MACRO block_546x675_107
   SIZE 207.48 BY 128.25 ;
END block_546x675_107

MACRO block_341x369_76
   SIZE 129.58 BY 70.11 ;
END block_341x369_76

MACRO block_414x1071_178
   SIZE 157.32 BY 203.49 ;
END block_414x1071_178

MACRO block_341x369_72
   SIZE 129.58 BY 70.11 ;
END block_341x369_72

MACRO block_535x747_102
   SIZE 203.3 BY 141.93 ;
END block_535x747_102

MACRO block_197x171_32
   SIZE 74.86 BY 32.49 ;
END block_197x171_32

MACRO block_671x747_104
   SIZE 254.98 BY 141.93 ;
END block_671x747_104

MACRO block_546x675_83
   SIZE 207.48 BY 128.25 ;
END block_546x675_83

MACRO block_197x171_33
   SIZE 74.86 BY 32.49 ;
END block_197x171_33

MACRO block_779x1125_90
   SIZE 296.02 BY 213.75 ;
END block_779x1125_90

MACRO block_159x2349_160
   SIZE 60.42 BY 446.31 ;
END block_159x2349_160

MACRO block_252x2349_162
   SIZE 95.76 BY 446.31 ;
END block_252x2349_162

MACRO block_348x2349_165
   SIZE 132.24 BY 446.31 ;
END block_348x2349_165

MACRO block_414x1917_342
   SIZE 157.32 BY 364.23 ;
END block_414x1917_342

MACRO block_546x675_77
   SIZE 207.48 BY 128.25 ;
END block_546x675_77

MACRO block_414x2007_358
   SIZE 157.32 BY 381.33 ;
END block_414x2007_358

MACRO block_546x675_97
   SIZE 207.48 BY 128.25 ;
END block_546x675_97

MACRO block_414x2007_358f
   SIZE 157.32 BY 381.33 ;
END block_414x2007_358f

MACRO block_575x801_42
   SIZE 218.5 BY 152.19 ;
END block_575x801_42

MACRO block_737x900_321
   SIZE 280.06 BY 171.0 ;
END block_737x900_321

MACRO block_644x675_89
   SIZE 244.72 BY 128.25 ;
END block_644x675_89

MACRO block_321x324_66
   SIZE 121.98 BY 61.56 ;
END block_321x324_66

MACRO block_567x774_60
   SIZE 215.46 BY 147.06 ;
END block_567x774_60

MACRO block_575x801_43
   SIZE 218.5 BY 152.19 ;
END block_575x801_43

MACRO block_567x774_62
   SIZE 215.46 BY 147.06 ;
END block_567x774_62

MACRO block_575x558_34
   SIZE 218.5 BY 106.02 ;
END block_575x558_34

MACRO block_126x2196_149
   SIZE 47.88 BY 417.24 ;
END block_126x2196_149

MACRO block_126x2196_148
   SIZE 47.88 BY 417.24 ;
END block_126x2196_148

MACRO block_575x315_26
   SIZE 218.5 BY 59.85 ;
END block_575x315_26

MACRO block_575x315_27
   SIZE 218.5 BY 59.85 ;
END block_575x315_27

MACRO block_414x1746_310
   SIZE 157.32 BY 331.74 ;
END block_414x1746_310

MACRO block_341x369_75
   SIZE 129.58 BY 70.11 ;
END block_341x369_75

MACRO block_533x1125_87
   SIZE 202.54 BY 213.75 ;
END block_533x1125_87

MACRO block_341x369_74
   SIZE 129.58 BY 70.11 ;
END block_341x369_74

MACRO block_535x747_102f
   SIZE 203.3 BY 141.93 ;
END block_535x747_102f

MACRO block_546x675_88
   SIZE 207.48 BY 128.25 ;
END block_546x675_88

MACRO block_1100x1125_93
   SIZE 418.0 BY 213.75 ;
END block_1100x1125_93

MACRO block_315x2349_162
   SIZE 119.7 BY 446.31 ;
END block_315x2349_162

MACRO block_737x1152_453
   SIZE 280.06 BY 218.88 ;
END block_737x1152_453

MACRO block_321x315_66
   SIZE 121.98 BY 59.85 ;
END block_321x315_66

MACRO block_737x1845_682
   SIZE 280.06 BY 350.55 ;
END block_737x1845_682

MACRO block_644x666_102
   SIZE 244.72 BY 126.54 ;
END block_644x666_102

MACRO block_535x801_109
   SIZE 203.3 BY 152.19 ;
END block_535x801_109

MACRO block_1338x6831_672
   SIZE 508.44 BY 1297.89 ;
END block_1338x6831_672

MACRO block_416x441_117
   SIZE 158.08 BY 83.79 ;
END block_416x441_117

MACRO block_535x945_130
   SIZE 203.3 BY 179.55 ;
END block_535x945_130

MACRO block_533x1125_122
   SIZE 202.54 BY 213.75 ;
END block_533x1125_122

MACRO block_546x675_102
   SIZE 207.48 BY 128.25 ;
END block_546x675_102

MACRO block_1829x2160_148
   SIZE 695.02 BY 410.4 ;
END block_1829x2160_148

MACRO block_1338x2160_145
   SIZE 508.44 BY 410.4 ;
END block_1338x2160_145

MACRO block_1829x2502_263
   SIZE 695.02 BY 475.38 ;
END block_1829x2502_263

MACRO block_1338x1773_192
   SIZE 508.44 BY 336.87 ;
END block_1338x1773_192

MACRO block_315x1863_130
   SIZE 119.7 BY 353.97 ;
END block_315x1863_130

MACRO block_414x2520_454
   SIZE 157.32 BY 478.8 ;
END block_414x2520_454

MACRO block_737x810_273
   SIZE 280.06 BY 153.9 ;
END block_737x810_273

MACRO block_779x1035_113
   SIZE 296.02 BY 196.65 ;
END block_779x1035_113

MACRO block_546x675_94
   SIZE 207.48 BY 128.25 ;
END block_546x675_94

MACRO block_315x558_44
   SIZE 119.7 BY 106.02 ;
END block_315x558_44

MACRO block_222x1926_135
   SIZE 84.36 BY 365.94 ;
END block_222x1926_135

MACRO block_222x1926_134
   SIZE 84.36 BY 365.94 ;
END block_222x1926_134

MACRO block_222x2349_162
   SIZE 84.36 BY 446.31 ;
END block_222x2349_162

MACRO block_73x72_14
   SIZE 27.74 BY 13.68 ;
END block_73x72_14

MACRO block_23x9_0
   SIZE 8.74 BY 1.71 ;
END block_23x9_0

MACRO block_73x72_15
   SIZE 27.74 BY 13.68 ;
END block_73x72_15

MACRO block_26x9_0
   SIZE 9.88 BY 1.71 ;
END block_26x9_0

MACRO block_100x144_0
   SIZE 38.0 BY 27.36 ;
END block_100x144_0

MACRO block_43x63_0
   SIZE 16.34 BY 11.97 ;
END block_43x63_0

END LIBRARY
