MACRO block_533x1215_91
   SIZE 202.54 BY 230.85 ;
END block_533x1215_91

MACRO block_546x675_88
   SIZE 207.48 BY 128.25 ;
END block_546x675_88

MACRO block_341x369_74
   SIZE 129.58 BY 70.11 ;
END block_341x369_74

MACRO block_535x945_130
   SIZE 203.3 BY 179.55 ;
END block_535x945_130

MACRO block_197x171_33
   SIZE 74.86 BY 32.49 ;
END block_197x171_33

MACRO block_7596x3465_370
   SIZE 2886.48 BY 658.35 ;
END block_7596x3465_370

MACRO block_646x2655_74
   SIZE 245.48 BY 504.45 ;
END block_646x2655_74

MACRO block_533x3717_657
   SIZE 202.54 BY 706.23 ;
END block_533x3717_657

MACRO block_416x441_105
   SIZE 158.08 BY 83.79 ;
END block_416x441_105

MACRO block_779x1467_106
   SIZE 296.02 BY 278.73 ;
END block_779x1467_106

MACRO block_341x369_76
   SIZE 129.58 BY 70.11 ;
END block_341x369_76

MACRO block_535x549_99
   SIZE 203.3 BY 104.31 ;
END block_535x549_99

MACRO block_197x171_32
   SIZE 74.86 BY 32.49 ;
END block_197x171_32

MACRO block_779x2844_174
   SIZE 296.02 BY 540.36 ;
END block_779x2844_174

MACRO block_341x369_80
   SIZE 129.58 BY 70.11 ;
END block_341x369_80

MACRO block_2456x1746_322
   SIZE 933.28 BY 331.74 ;
END block_2456x1746_322

MACRO block_546x675_83
   SIZE 207.48 BY 128.25 ;
END block_546x675_83

MACRO block_341x369_84
   SIZE 129.58 BY 70.11 ;
END block_341x369_84

MACRO block_1657x2799_1266
   SIZE 629.66 BY 531.81 ;
END block_1657x2799_1266

MACRO block_644x666_91
   SIZE 244.72 BY 126.54 ;
END block_644x666_91

MACRO block_336x333_85
   SIZE 127.68 BY 63.27 ;
END block_336x333_85

MACRO block_414x1665_290
   SIZE 157.32 BY 316.35 ;
END block_414x1665_290

MACRO block_546x675_72
   SIZE 207.48 BY 128.25 ;
END block_546x675_72

MACRO block_341x369_71
   SIZE 129.58 BY 70.11 ;
END block_341x369_71

MACRO block_535x549_106
   SIZE 203.3 BY 104.31 ;
END block_535x549_106

MACRO block_779x5265_948
   SIZE 296.02 BY 1000.35 ;
END block_779x5265_948

MACRO block_416x441_108
   SIZE 158.08 BY 83.79 ;
END block_416x441_108

MACRO block_533x1125_122
   SIZE 202.54 BY 213.75 ;
END block_533x1125_122

MACRO block_1596x3978_542
   SIZE 606.48 BY 755.82 ;
END block_1596x3978_542

MACRO block_716x810_89
   SIZE 272.08 BY 153.9 ;
END block_716x810_89

MACRO block_232x297_54
   SIZE 88.16 BY 56.43 ;
END block_232x297_54

MACRO block_1338x1746_319
   SIZE 508.44 BY 331.74 ;
END block_1338x1746_319

MACRO block_546x675_87
   SIZE 207.48 BY 128.25 ;
END block_546x675_87

MACRO block_341x369_82
   SIZE 129.58 BY 70.11 ;
END block_341x369_82

MACRO block_1338x1746_319f
   SIZE 508.44 BY 331.74 ;
END block_1338x1746_319f

MACRO block_546x675_82
   SIZE 207.48 BY 128.25 ;
END block_546x675_82

MACRO block_2456x1746_322f
   SIZE 933.28 BY 331.74 ;
END block_2456x1746_322f

MACRO block_2456x1755_322
   SIZE 933.28 BY 333.45 ;
END block_2456x1755_322

MACRO block_546x675_77
   SIZE 207.48 BY 128.25 ;
END block_546x675_77

MACRO block_2456x6183_356
   SIZE 933.28 BY 1174.77 ;
END block_2456x6183_356

MACRO block_416x441_120
   SIZE 158.08 BY 83.79 ;
END block_416x441_120

MACRO block_2456x6183_356f
   SIZE 933.28 BY 1174.77 ;
END block_2456x6183_356f

MACRO block_779x1125_90
   SIZE 296.02 BY 213.75 ;
END block_779x1125_90

MACRO block_535x747_156
   SIZE 203.3 BY 141.93 ;
END block_535x747_156

MACRO block_546x675_78
   SIZE 207.48 BY 128.25 ;
END block_546x675_78

MACRO block_2953x3276_1641
   SIZE 1122.14 BY 622.44 ;
END block_2953x3276_1641

MACRO block_644x666_92
   SIZE 244.72 BY 126.54 ;
END block_644x666_92

MACRO block_336x333_86
   SIZE 127.68 BY 63.27 ;
END block_336x333_86

MACRO block_414x1962_350
   SIZE 157.32 BY 372.78 ;
END block_414x1962_350

MACRO block_546x675_73
   SIZE 207.48 BY 128.25 ;
END block_546x675_73

MACRO block_126x2403_162
   SIZE 47.88 BY 456.57 ;
END block_126x2403_162

MACRO block_3369x4428_2245
   SIZE 1280.22 BY 841.32 ;
END block_3369x4428_2245

MACRO block_345x378_86
   SIZE 131.1 BY 71.82 ;
END block_345x378_86

MACRO block_779x5571_1004
   SIZE 296.02 BY 1058.49 ;
END block_779x5571_1004

MACRO block_416x432_108
   SIZE 158.08 BY 82.08 ;
END block_416x432_108

MACRO block_779x5571_1004f
   SIZE 296.02 BY 1058.49 ;
END block_779x5571_1004f

MACRO block_189x1980_137
   SIZE 71.82 BY 376.2 ;
END block_189x1980_137

MACRO block_189x1980_136
   SIZE 71.82 BY 376.2 ;
END block_189x1980_136

MACRO block_533x1188_205
   SIZE 202.54 BY 225.72 ;
END block_533x1188_205

MACRO block_779x1296_98
   SIZE 296.02 BY 246.24 ;
END block_779x1296_98

MACRO block_1338x1683_180
   SIZE 508.44 BY 319.77 ;
END block_1338x1683_180

MACRO block_341x369_77
   SIZE 129.58 BY 70.11 ;
END block_341x369_77

MACRO block_779x1386_102
   SIZE 296.02 BY 263.34 ;
END block_779x1386_102

MACRO block_414x1620_282
   SIZE 157.32 BY 307.8 ;
END block_414x1620_282

MACRO block_341x369_72
   SIZE 129.58 BY 70.11 ;
END block_341x369_72

MACRO block_575x441_31
   SIZE 218.5 BY 83.79 ;
END block_575x441_31

MACRO block_414x4230_750
   SIZE 157.32 BY 803.7 ;
END block_414x4230_750

MACRO block_416x441_104
   SIZE 158.08 BY 83.79 ;
END block_416x441_104

MACRO block_414x1701_298
   SIZE 157.32 BY 323.19 ;
END block_414x1701_298

MACRO block_126x2043_138
   SIZE 47.88 BY 388.17 ;
END block_126x2043_138

MACRO block_414x1431_246
   SIZE 157.32 BY 271.89 ;
END block_414x1431_246

MACRO block_414x1431_246f
   SIZE 157.32 BY 271.89 ;
END block_414x1431_246f

MACRO block_1591x2133_394
   SIZE 604.58 BY 405.27 ;
END block_1591x2133_394

MACRO block_1338x1773_192
   SIZE 508.44 BY 336.87 ;
END block_1338x1773_192

MACRO block_1009x918_401
   SIZE 383.42 BY 174.42 ;
END block_1009x918_401

MACRO block_644x666_90
   SIZE 244.72 BY 126.54 ;
END block_644x666_90

MACRO block_294x270_66
   SIZE 111.72 BY 51.3 ;
END block_294x270_66

MACRO block_323x801_41
   SIZE 122.74 BY 152.19 ;
END block_323x801_41

MACRO block_126x1863_126
   SIZE 47.88 BY 353.97 ;
END block_126x1863_126

MACRO block_535x846_184
   SIZE 203.3 BY 160.74 ;
END block_535x846_184

MACRO block_414x1035_170
   SIZE 157.32 BY 196.65 ;
END block_414x1035_170

MACRO block_341x369_68
   SIZE 129.58 BY 70.11 ;
END block_341x369_68

MACRO block_126x1080_74
   SIZE 47.88 BY 205.2 ;
END block_126x1080_74

MACRO block_414x2565_462
   SIZE 157.32 BY 487.35 ;
END block_414x2565_462

MACRO block_341x369_75
   SIZE 129.58 BY 70.11 ;
END block_341x369_75

MACRO block_414x5220_934
   SIZE 157.32 BY 991.8 ;
END block_414x5220_934

MACRO block_189x2259_154
   SIZE 71.82 BY 429.21 ;
END block_189x2259_154

MACRO block_189x2313_158
   SIZE 71.82 BY 439.47 ;
END block_189x2313_158

MACRO block_414x6129_1110
   SIZE 157.32 BY 1164.51 ;
END block_414x6129_1110

MACRO block_416x441_112
   SIZE 158.08 BY 83.79 ;
END block_416x441_112

MACRO block_414x6129_1110f
   SIZE 157.32 BY 1164.51 ;
END block_414x6129_1110f

MACRO block_126x1710_116
   SIZE 47.88 BY 324.9 ;
END block_126x1710_116

MACRO block_535x801_170
   SIZE 203.3 BY 152.19 ;
END block_535x801_170

MACRO block_414x3519_618
   SIZE 157.32 BY 668.61 ;
END block_414x3519_618

MACRO block_414x3519_618f
   SIZE 157.32 BY 668.61 ;
END block_414x3519_618f

MACRO block_1004x3474_655
   SIZE 381.52 BY 660.06 ;
END block_1004x3474_655

MACRO block_1004x3474_656
   SIZE 381.52 BY 660.06 ;
END block_1004x3474_656

MACRO block_73x72_14
   SIZE 27.74 BY 13.68 ;
END block_73x72_14

END LIBRARY
