MACRO block_4449x4239_2703
   SIZE 1690.62 BY 805.41 ;
END block_4449x4239_2703

MACRO block_423x405_126
   SIZE 160.74 BY 76.95 ;
END block_423x405_126

MACRO block_644x666_97
   SIZE 244.72 BY 126.54 ;
END block_644x666_97

MACRO block_1100x1746_319
   SIZE 418.0 BY 331.74 ;
END block_1100x1746_319

MACRO block_546x675_72
   SIZE 207.48 BY 128.25 ;
END block_546x675_72

MACRO block_341x369_81
   SIZE 129.58 BY 70.11 ;
END block_341x369_81

MACRO block_341x369_82
   SIZE 129.58 BY 70.11 ;
END block_341x369_82

MACRO block_1100x1746_319f
   SIZE 418.0 BY 331.74 ;
END block_1100x1746_319f

MACRO block_546x675_77
   SIZE 207.48 BY 128.25 ;
END block_546x675_77

MACRO block_546x675_73
   SIZE 207.48 BY 128.25 ;
END block_546x675_73

MACRO block_2953x4239_2403
   SIZE 1122.14 BY 805.41 ;
END block_2953x4239_2403

MACRO block_336x333_86
   SIZE 127.68 BY 63.27 ;
END block_336x333_86

MACRO block_533x1080_118
   SIZE 202.54 BY 205.2 ;
END block_533x1080_118

MACRO block_341x369_74
   SIZE 129.58 BY 70.11 ;
END block_341x369_74

MACRO block_546x675_108
   SIZE 207.48 BY 128.25 ;
END block_546x675_108

MACRO block_644x666_98
   SIZE 244.72 BY 126.54 ;
END block_644x666_98

MACRO block_533x1080_118f
   SIZE 202.54 BY 205.2 ;
END block_533x1080_118f

MACRO block_341x369_73
   SIZE 129.58 BY 70.11 ;
END block_341x369_73

MACRO block_73x72_14
   SIZE 27.74 BY 13.68 ;
END block_73x72_14

MACRO block_73x72_15
   SIZE 27.74 BY 13.68 ;
END block_73x72_15

END LIBRARY
