MACRO MAS4439
     SIZE 53.300 BY 196.200 ;
END MAS4439

MACRO MAS4440
     SIZE 54.600 BY 67.500 ;
END MAS4440

MACRO MAS4441
     SIZE 34.100 BY 36.900 ;
END MAS4441

MACRO MAS4447
     SIZE 32.300 BY 44.100 ;
END MAS4447

MACRO MAS4448
     SIZE 53.300 BY 134.100 ;
END MAS4448

MACRO MAS4449
     SIZE 34.100 BY 36.900 ;
END MAS4449

MACRO MAS4453
     SIZE 73.700 BY 90.900 ;
END MAS4453

MACRO MAS4454
     SIZE 64.400 BY 66.600 ;
END MAS4454

MACRO MAS4455
     SIZE 32.100 BY 32.400 ;
END MAS4455

MACRO MAS4457
     SIZE 31.500 BY 144.000 ;
END MAS4457

MACRO MAS4459
     SIZE 100.900 BY 90.900 ;
END MAS4459

MACRO MAS4460
     SIZE 64.400 BY 66.600 ;
END MAS4460

MACRO MAS4461
     SIZE 29.400 BY 27.000 ;
END MAS4461

MACRO MAS4463
     SIZE 73.700 BY 90.900 ;
END MAS4463

MACRO MAS4464
     SIZE 32.100 BY 32.400 ;
END MAS4464

MACRO MAS4466
     SIZE 100.900 BY 90.900 ;
END MAS4466

MACRO MAS4467
     SIZE 29.400 BY 27.000 ;
END MAS4467

MACRO MAS4469
     SIZE 100.900 BY 90.000 ;
END MAS4469

MACRO MAS4470
     SIZE 64.400 BY 67.500 ;
END MAS4470

MACRO MAS4471
     SIZE 29.400 BY 27.900 ;
END MAS4471

MACRO MAS4472
     SIZE 73.700 BY 90.000 ;
END MAS4472

MACRO MAS4473
     SIZE 32.100 BY 31.500 ;
END MAS4473

MACRO MAS4474
     SIZE 100.900 BY 90.000 ;
END MAS4474

MACRO MAS4476
     SIZE 100.900 BY 90.000 ;
END MAS4476

MACRO MAS4477
     SIZE 73.700 BY 90.000 ;
END MAS4477

MACRO MAS4478
     SIZE 32.100 BY 31.500 ;
END MAS4478

MACRO MAS4479
     SIZE 100.900 BY 90.000 ;
END MAS4479

MACRO MAS4483
     SIZE 31.500 BY 243.900 ;
END MAS4483

MACRO MAS4484
     SIZE 31.500 BY 243.900 ;
END MAS4484

MACRO MAS4489
     SIZE 87.600 BY 387.900 ;
END MAS4489

MACRO MAS4490
     SIZE 54.600 BY 67.500 ;
END MAS4490

MACRO MAS4491
     SIZE 23.200 BY 29.700 ;
END MAS4491

MACRO MAS4492
     SIZE 87.600 BY 387.900 ;
END MAS4492

MACRO MAS4493
     SIZE 23.200 BY 29.700 ;
END MAS4493

MACRO MAS4494
     SIZE 87.600 BY 388.800 ;
END MAS4494

MACRO MAS4495
     SIZE 23.200 BY 29.700 ;
END MAS4495

MACRO MAS4496
     SIZE 87.600 BY 387.000 ;
END MAS4496

MACRO MAS4497
     SIZE 87.600 BY 387.900 ;
END MAS4497

MACRO MAS4498
     SIZE 87.600 BY 387.900 ;
END MAS4498

MACRO MAS4499
     SIZE 23.200 BY 29.700 ;
END MAS4499

MACRO MAS4500
     SIZE 87.600 BY 388.800 ;
END MAS4500

MACRO MAS4501
     SIZE 87.600 BY 388.800 ;
END MAS4501

MACRO MAS4502
     SIZE 41.200 BY 765.900 ;
END MAS4502

MACRO MAS4503
     SIZE 71.600 BY 81.000 ;
END MAS4503

MACRO MAS4504
     SIZE 29.200 BY 35.100 ;
END MAS4504

MACRO MAS4505
     SIZE 41.200 BY 765.000 ;
END MAS4505

MACRO MAS4506
     SIZE 29.200 BY 36.000 ;
END MAS4506

MACRO MAS4507
     SIZE 41.200 BY 765.000 ;
END MAS4507

MACRO MAS4508
     SIZE 41.200 BY 765.000 ;
END MAS4508

MACRO MAS4509
     SIZE 29.200 BY 36.000 ;
END MAS4509

MACRO MAS4510
     SIZE 41.200 BY 765.000 ;
END MAS4510

MACRO MAS4511
     SIZE 29.200 BY 36.000 ;
END MAS4511

MACRO MAS4512
     SIZE 41.200 BY 765.000 ;
END MAS4512

MACRO MAS4514
     SIZE 18.900 BY 259.200 ;
END MAS4514

MACRO MAS4515
     SIZE 18.900 BY 259.200 ;
END MAS4515

MACRO MAS4516
     SIZE 18.900 BY 110.700 ;
END MAS4516

MACRO MAS4518
     SIZE 31.500 BY 119.700 ;
END MAS4518

MACRO MAS4520
     SIZE 31.500 BY 119.700 ;
END MAS4520

MACRO MAS4521
     SIZE 18.900 BY 252.900 ;
END MAS4521

MACRO MAS4523
     SIZE 18.900 BY 252.900 ;
END MAS4523

MACRO MAS4524
     SIZE 31.500 BY 173.700 ;
END MAS4524

MACRO MAS4525
     SIZE 31.500 BY 173.700 ;
END MAS4525

MACRO MAS4526
     SIZE 18.900 BY 110.700 ;
END MAS4526

MACRO MAS4527
     SIZE 31.500 BY 119.700 ;
END MAS4527

MACRO MAS4528
     SIZE 29.400 BY 27.000 ;
END MAS4528

MACRO MAS4529
     SIZE 73.700 BY 90.900 ;
END MAS4529

MACRO MAS4530
     SIZE 32.100 BY 32.400 ;
END MAS4530

MACRO MAS4532
     SIZE 29.400 BY 27.000 ;
END MAS4532

MACRO MAS4533
     SIZE 64.400 BY 66.600 ;
END MAS4533

MACRO MAS4534
     SIZE 73.700 BY 90.000 ;
END MAS4534

MACRO MAS4535
     SIZE 12.600 BY 92.700 ;
END MAS4535

MACRO MAS4536
     SIZE 31.500 BY 173.700 ;
END MAS4536

MACRO MAS4537
     SIZE 40.400 BY 208.800 ;
END MAS4537

MACRO MAS4538
     SIZE 71.600 BY 81.000 ;
END MAS4538

MACRO MAS4539
     SIZE 21.700 BY 20.700 ;
END MAS4539

MACRO MAS4540
     SIZE 40.400 BY 778.500 ;
END MAS4540

MACRO MAS4541
     SIZE 29.200 BY 35.100 ;
END MAS4541

MACRO MAS4542
     SIZE 18.900 BY 110.700 ;
END MAS4542

MACRO MAS4543
     SIZE 31.500 BY 119.700 ;
END MAS4543

MACRO MAS4544
     SIZE 18.900 BY 252.900 ;
END MAS4544

MACRO MAS4545
     SIZE 12.600 BY 237.600 ;
END MAS4545

MACRO MAS4546
     SIZE 12.600 BY 237.600 ;
END MAS4546

MACRO MAS4547
     SIZE 12.600 BY 237.600 ;
END MAS4547

MACRO MAS4572
     SIZE 7.300 BY 7.200 ;
END MAS4572

MACRO MAS4718
     SIZE 7.300 BY 7.200 ;
END MAS4718

END LIBRARY
