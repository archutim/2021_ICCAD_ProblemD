MACRO block_414x2007_358
   SIZE 157.32 BY 381.33 ;
END block_414x2007_358

MACRO block_341x369_76
   SIZE 129.58 BY 70.11 ;
END block_341x369_76

MACRO block_737x1845_682
   SIZE 280.06 BY 350.55 ;
END block_737x1845_682

MACRO block_644x666_92
   SIZE 244.72 BY 126.54 ;
END block_644x666_92

MACRO block_321x315_66
   SIZE 121.98 BY 59.85 ;
END block_321x315_66

MACRO block_779x1431_153
   SIZE 296.02 BY 271.89 ;
END block_779x1431_153

MACRO block_546x675_104
   SIZE 207.48 BY 128.25 ;
END block_546x675_104

MACRO block_533x1044_173
   SIZE 202.54 BY 198.36 ;
END block_533x1044_173

MACRO block_341x369_70
   SIZE 129.58 BY 70.11 ;
END block_341x369_70

MACRO block_779x2502_158
   SIZE 296.02 BY 475.38 ;
END block_779x2502_158

MACRO block_341x369_80
   SIZE 129.58 BY 70.11 ;
END block_341x369_80

MACRO block_1024x2502_161
   SIZE 389.12 BY 475.38 ;
END block_1024x2502_161

MACRO block_341x369_82
   SIZE 129.58 BY 70.11 ;
END block_341x369_82

MACRO block_414x1746_310
   SIZE 157.32 BY 331.74 ;
END block_414x1746_310

MACRO block_341x369_75
   SIZE 129.58 BY 70.11 ;
END block_341x369_75

MACRO block_533x1125_87
   SIZE 202.54 BY 213.75 ;
END block_533x1125_87

MACRO block_341x369_74
   SIZE 129.58 BY 70.11 ;
END block_341x369_74

MACRO block_126x648_46
   SIZE 47.88 BY 123.12 ;
END block_126x648_46

MACRO block_535x945_130
   SIZE 203.3 BY 179.55 ;
END block_535x945_130

MACRO block_546x675_105
   SIZE 207.48 BY 128.25 ;
END block_546x675_105

MACRO block_197x171_33
   SIZE 74.86 BY 32.49 ;
END block_197x171_33

MACRO block_2456x4626_834
   SIZE 933.28 BY 878.94 ;
END block_2456x4626_834

MACRO block_416x441_112
   SIZE 158.08 BY 83.79 ;
END block_416x441_112

MACRO block_126x351_27
   SIZE 47.88 BY 66.69 ;
END block_126x351_27

MACRO block_533x1539_269
   SIZE 202.54 BY 292.41 ;
END block_533x1539_269

MACRO block_671x801_111
   SIZE 254.98 BY 152.19 ;
END block_671x801_111

MACRO block_197x180_33
   SIZE 74.86 BY 34.2 ;
END block_197x180_33

MACRO block_1338x2160_145
   SIZE 508.44 BY 410.4 ;
END block_1338x2160_145

MACRO block_533x1125_122
   SIZE 202.54 BY 213.75 ;
END block_533x1125_122

MACRO block_1829x2160_148
   SIZE 695.02 BY 410.4 ;
END block_1829x2160_148

MACRO block_341x369_84
   SIZE 129.58 BY 70.11 ;
END block_341x369_84

MACRO block_779x1467_106
   SIZE 296.02 BY 278.73 ;
END block_779x1467_106

MACRO block_1829x2502_263
   SIZE 695.02 BY 475.38 ;
END block_1829x2502_263

MACRO block_1338x1773_192
   SIZE 508.44 BY 336.87 ;
END block_1338x1773_192

MACRO block_546x684_100
   SIZE 207.48 BY 129.96 ;
END block_546x684_100

MACRO block_737x1152_453
   SIZE 280.06 BY 218.88 ;
END block_737x1152_453

MACRO block_644x666_91
   SIZE 244.72 BY 126.54 ;
END block_644x666_91

MACRO block_321x324_66
   SIZE 121.98 BY 61.56 ;
END block_321x324_66

MACRO block_315x1863_130
   SIZE 119.7 BY 353.97 ;
END block_315x1863_130

MACRO block_96x2070_138
   SIZE 36.48 BY 393.3 ;
END block_96x2070_138

MACRO block_737x3078_1192
   SIZE 280.06 BY 584.82 ;
END block_737x3078_1192

MACRO block_644x675_93
   SIZE 244.72 BY 128.25 ;
END block_644x675_93

MACRO block_321x324_65
   SIZE 121.98 BY 61.56 ;
END block_321x324_65

MACRO block_779x1557_110
   SIZE 296.02 BY 295.83 ;
END block_779x1557_110

MACRO block_315x558_44
   SIZE 119.7 BY 106.02 ;
END block_315x558_44

MACRO block_414x3978_702
   SIZE 157.32 BY 755.82 ;
END block_414x3978_702

MACRO block_416x441_104
   SIZE 158.08 BY 83.79 ;
END block_416x441_104

MACRO block_414x3969_702
   SIZE 157.32 BY 754.11 ;
 END block_414x3969_702

MACRO block_737x819_279
   SIZE 280.06 BY 155.61 ;
END block_737x819_279

MACRO block_1100x1557_168
   SIZE 418.0 BY 295.83 ;
END block_1100x1557_168

MACRO block_341x369_78
   SIZE 129.58 BY 70.11 ;
END block_341x369_78

MACRO block_315x981_72
   SIZE 119.7 BY 186.39 ;
END block_315x981_72

MACRO block_535x756_102
   SIZE 203.3 BY 143.64 ;
END block_535x756_102

MACRO block_197x180_32
   SIZE 74.86 BY 34.2 ;
END block_197x180_32

MACRO block_533x4428_789
   SIZE 202.54 BY 841.32 ;
END block_533x4428_789

MACRO block_533x4428_789f
   SIZE 202.54 BY 841.32 ;
END block_533x4428_789f

MACRO block_416x450_106
   SIZE 158.08 BY 85.5 ;
END block_416x450_106

MACRO block_416x441_106
   SIZE 158.08 BY 83.79 ;
END block_416x441_106

MACRO block_315x2106_146
   SIZE 119.7 BY 400.14 ;
END block_315x2106_146

MACRO block_73x72_14
   SIZE 27.74 BY 13.68 ;
END block_73x72_14

MACRO block_73x72_15
   SIZE 27.74 BY 13.68 ;
END block_73x72_15

END LIBRARY
