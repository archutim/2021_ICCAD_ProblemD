MACRO MAS4584
     SIZE 230.500 BY 90.000 ;
END MAS4584

MACRO MAS4585
     SIZE 33.600 BY 33.300 ;
END MAS4585

MACRO MAS4586
     SIZE 230.500 BY 90.000 ;
END MAS4586

MACRO MAS4587
     SIZE 64.400 BY 66.600 ;
END MAS4587

MACRO MAS4588
     SIZE 33.600 BY 33.300 ;
END MAS4588

MACRO MAS4589
     SIZE 230.500 BY 90.000 ;
END MAS4589

MACRO MAS4590
     SIZE 64.400 BY 66.600 ;
END MAS4590

MACRO MAS4591
     SIZE 64.400 BY 66.600 ;
END MAS4591

MACRO MAS4592
     SIZE 33.600 BY 33.300 ;
END MAS4592

MACRO MAS4593
     SIZE 33.600 BY 33.300 ;
END MAS4593

MACRO MAS4594
     SIZE 230.500 BY 90.000 ;
END MAS4594

MACRO MAS4595
     SIZE 64.400 BY 66.600 ;
END MAS4595

MACRO MAS4596
     SIZE 33.600 BY 33.300 ;
END MAS4596

MACRO MAS4597
     SIZE 33.600 BY 32.400 ;
END MAS4597

MACRO MAS4598
     SIZE 64.400 BY 66.600 ;
END MAS4598

MACRO MAS4599
     SIZE 33.600 BY 33.300 ;
END MAS4599

MACRO MAS4600
     SIZE 230.500 BY 89.100 ;
END MAS4600

MACRO MAS4601
     SIZE 64.400 BY 67.500 ;
END MAS4601

MACRO MAS4602
     SIZE 230.500 BY 90.000 ;
END MAS4602

MACRO MAS4603
     SIZE 64.400 BY 67.500 ;
END MAS4603

MACRO MAS4604
     SIZE 44.100 BY 92.700 ;
END MAS4604

MACRO MAS4605
     SIZE 45.200 BY 774.900 ;
END MAS4605

MACRO MAS4606
     SIZE 71.600 BY 81.000 ;
END MAS4606

MACRO MAS4607
     SIZE 29.200 BY 34.200 ;
END MAS4607

MACRO MAS4608
     SIZE 45.200 BY 774.900 ;
END MAS4608

MACRO MAS4609
     SIZE 29.200 BY 36.000 ;
END MAS4609

MACRO MAS4610
     SIZE 42.000 BY 760.500 ;
END MAS4610

MACRO MAS4611
     SIZE 29.200 BY 35.100 ;
END MAS4611

MACRO MAS4612
     SIZE 42.000 BY 760.500 ;
END MAS4612

MACRO MAS4613
     SIZE 29.200 BY 36.000 ;
END MAS4613

MACRO MAS4614
     SIZE 42.000 BY 760.500 ;
END MAS4614

MACRO MAS4615
     SIZE 71.600 BY 81.000 ;
END MAS4615

MACRO MAS4616
     SIZE 29.200 BY 35.100 ;
END MAS4616

MACRO MAS4617
     SIZE 42.000 BY 760.500 ;
END MAS4617

MACRO MAS4618
     SIZE 29.200 BY 35.100 ;
END MAS4618

MACRO MAS4619
     SIZE 42.000 BY 760.500 ;
END MAS4619

MACRO MAS4620
     SIZE 42.000 BY 760.500 ;
END MAS4620

MACRO MAS4621
     SIZE 29.200 BY 35.100 ;
END MAS4621

MACRO MAS4622
     SIZE 42.000 BY 760.500 ;
END MAS4622

MACRO MAS4623
     SIZE 29.200 BY 35.100 ;
END MAS4623

MACRO MAS4624
     SIZE 42.000 BY 760.500 ;
END MAS4624

MACRO MAS4625
     SIZE 29.200 BY 35.100 ;
END MAS4625

MACRO MAS4626
     SIZE 44.100 BY 213.300 ;
END MAS4626

MACRO MAS4627
     SIZE 44.100 BY 213.300 ;
END MAS4627

MACRO MAS4628
     SIZE 31.500 BY 92.700 ;
END MAS4628

MACRO MAS4629
     SIZE 44.100 BY 104.400 ;
END MAS4629

MACRO MAS4630
     SIZE 7.300 BY 7.200 ;
END MAS4630

MACRO MAS4631
     SIZE 7.300 BY 7.200 ;
END MAS4631

END LIBRARY
