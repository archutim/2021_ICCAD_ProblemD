MACRO MAS4478
     SIZE 47.400 BY 599.400 ;
END MAS4478

MACRO MAS4479
     SIZE 54.600 BY 68.400 ;
END MAS4479

MACRO MAS4480
     SIZE 41.600 BY 44.100 ;
END MAS4480

MACRO MAS4481
     SIZE 557.200 BY 612.900 ;
END MAS4481

MACRO MAS4482
     SIZE 64.600 BY 265.500 ;
END MAS4482

MACRO MAS4483
     SIZE 53.300 BY 337.500 ;
END MAS4483

MACRO MAS4484
     SIZE 41.600 BY 44.100 ;
END MAS4484

MACRO MAS4485
     SIZE 108.400 BY 340.200 ;
END MAS4485

MACRO MAS4486
     SIZE 23.200 BY 29.700 ;
END MAS4486

MACRO MAS4487
     SIZE 108.400 BY 263.700 ;
END MAS4487

MACRO MAS4488
     SIZE 71.600 BY 81.900 ;
END MAS4488

MACRO MAS4489
     SIZE 23.200 BY 29.700 ;
END MAS4489

MACRO MAS4490
     SIZE 58.800 BY 204.300 ;
END MAS4490

MACRO MAS4491
     SIZE 71.600 BY 81.900 ;
END MAS4491

MACRO MAS4492
     SIZE 21.700 BY 20.700 ;
END MAS4492

MACRO MAS4493
     SIZE 38.900 BY 118.800 ;
END MAS4493

MACRO MAS4494
     SIZE 77.900 BY 177.300 ;
END MAS4494

MACRO MAS4495
     SIZE 34.100 BY 36.900 ;
END MAS4495

MACRO MAS4496
     SIZE 58.800 BY 194.400 ;
END MAS4496

MACRO MAS4497
     SIZE 71.600 BY 81.000 ;
END MAS4497

MACRO MAS4498
     SIZE 21.700 BY 20.700 ;
END MAS4498

MACRO MAS4499
     SIZE 77.900 BY 171.000 ;
END MAS4499

MACRO MAS4500
     SIZE 54.600 BY 68.400 ;
END MAS4500

MACRO MAS4501
     SIZE 34.100 BY 36.000 ;
END MAS4501

MACRO MAS4502
     SIZE 58.800 BY 195.300 ;
END MAS4502

MACRO MAS4503
     SIZE 21.700 BY 21.600 ;
END MAS4503

MACRO MAS4504
     SIZE 230.500 BY 301.500 ;
END MAS4504

MACRO MAS4505
     SIZE 64.400 BY 67.500 ;
END MAS4505

MACRO MAS4506
     SIZE 33.600 BY 33.300 ;
END MAS4506

MACRO MAS4507
     SIZE 230.500 BY 301.500 ;
END MAS4507

MACRO MAS4508
     SIZE 33.600 BY 33.300 ;
END MAS4508

MACRO MAS4509
     SIZE 49.200 BY 117.900 ;
END MAS4509

MACRO MAS4510
     SIZE 19.700 BY 18.000 ;
END MAS4510

MACRO MAS4511
     SIZE 58.800 BY 112.500 ;
END MAS4511

MACRO MAS4512
     SIZE 19.700 BY 17.100 ;
END MAS4512

MACRO MAS4513
     SIZE 49.200 BY 131.400 ;
END MAS4513

MACRO MAS4514
     SIZE 19.700 BY 17.100 ;
END MAS4514

MACRO MAS4515
     SIZE 77.900 BY 610.200 ;
END MAS4515

MACRO MAS4516
     SIZE 41.600 BY 44.100 ;
END MAS4516

MACRO MAS4517
     SIZE 77.900 BY 610.200 ;
END MAS4517

MACRO MAS4518
     SIZE 77.900 BY 610.200 ;
END MAS4518

MACRO MAS4519
     SIZE 77.900 BY 610.200 ;
END MAS4519

MACRO MAS4520
     SIZE 54.600 BY 68.400 ;
END MAS4520

MACRO MAS4521
     SIZE 41.600 BY 44.100 ;
END MAS4521

MACRO MAS4522
     SIZE 77.900 BY 610.200 ;
END MAS4522

MACRO MAS4523
     SIZE 41.600 BY 43.200 ;
END MAS4523

MACRO MAS4524
     SIZE 77.900 BY 610.200 ;
END MAS4524

MACRO MAS4525
     SIZE 77.900 BY 610.200 ;
END MAS4525

MACRO MAS4526
     SIZE 77.900 BY 610.200 ;
END MAS4526

MACRO MAS4527
     SIZE 54.600 BY 67.500 ;
END MAS4527

MACRO MAS4528
     SIZE 49.200 BY 122.400 ;
END MAS4528

MACRO MAS4529
     SIZE 71.600 BY 81.900 ;
END MAS4529

MACRO MAS4530
     SIZE 19.700 BY 18.000 ;
END MAS4530

MACRO MAS4531
     SIZE 12.600 BY 189.000 ;
END MAS4531

MACRO MAS4532
     SIZE 18.900 BY 225.900 ;
END MAS4532

MACRO MAS4533
     SIZE 18.900 BY 225.900 ;
END MAS4533

MACRO MAS4534
     SIZE 18.900 BY 210.600 ;
END MAS4534

MACRO MAS4535
     SIZE 18.900 BY 210.600 ;
END MAS4535

MACRO MAS4536
     SIZE 12.600 BY 177.300 ;
END MAS4536

MACRO MAS4537
     SIZE 12.600 BY 55.800 ;
END MAS4537

MACRO MAS4538
     SIZE 12.600 BY 146.700 ;
END MAS4538

MACRO MAS4539
     SIZE 18.900 BY 255.600 ;
END MAS4539

MACRO MAS4540
     SIZE 18.900 BY 255.600 ;
END MAS4540

MACRO MAS4541
     SIZE 18.900 BY 246.600 ;
END MAS4541

MACRO MAS4542
     SIZE 18.900 BY 246.600 ;
END MAS4542

MACRO MAS4543
     SIZE 7.300 BY 7.200 ;
END MAS4543

MACRO MAS4544
     SIZE 7.300 BY 7.200 ;
END MAS4544

END LIBRARY
