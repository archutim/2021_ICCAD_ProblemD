MACRO MAS1901
     SIZE 37.800 BY 210.600 ;
END MAS1901

MACRO MAS1902
     SIZE 37.800 BY 210.600 ;
END MAS1902

MACRO MAS1903
     SIZE 37.800 BY 225.900 ;
END MAS1903

MACRO MAS1904
     SIZE 370.000 BY 612.900 ;
END MAS1904

MACRO MAS1905
     SIZE 64.600 BY 266.400 ;
END MAS1905

MACRO MAS1906
     SIZE 56.700 BY 59.400 ;
END MAS1906

MACRO MAS1907
     SIZE 37.800 BY 210.600 ;
END MAS1907

MACRO MAS1908
     SIZE 37.800 BY 216.900 ;
END MAS1908

MACRO MAS1909
     SIZE 37.800 BY 216.900 ;
END MAS1909

MACRO MAS1910
     SIZE 12.600 BY 210.600 ;
END MAS1910

MACRO MAS1911
     SIZE 12.600 BY 210.600 ;
END MAS1911

MACRO MAS1912
     SIZE 18.900 BY 113.400 ;
END MAS1912

MACRO MAS1913
     SIZE 22.200 BY 210.600 ;
END MAS1913

MACRO MAS1914
     SIZE 245.600 BY 280.800 ;
END MAS1914

MACRO MAS1915
     SIZE 54.600 BY 68.400 ;
END MAS1915

MACRO MAS1916
     SIZE 34.100 BY 36.900 ;
END MAS1916

MACRO MAS1917
     SIZE 54.600 BY 68.400 ;
END MAS1917

MACRO MAS1918
     SIZE 22.200 BY 210.600 ;
END MAS1918

MACRO MAS1919
     SIZE 18.900 BY 113.400 ;
END MAS1919

MACRO MAS1920
     SIZE 77.900 BY 265.500 ;
END MAS1920

MACRO MAS1921
     SIZE 77.900 BY 265.500 ;
END MAS1921

MACRO MAS1922
     SIZE 77.900 BY 265.500 ;
END MAS1922

MACRO MAS1924
     SIZE 34.100 BY 36.900 ;
END MAS1924

MACRO MAS1925
     SIZE 34.100 BY 36.900 ;
END MAS1925

MACRO MAS1926
     SIZE 29.200 BY 36.000 ;
END MAS1926

MACRO MAS1927
     SIZE 71.600 BY 81.900 ;
END MAS1927

MACRO MAS1928
     SIZE 53.200 BY 765.000 ;
END MAS1928

MACRO MAS1929
     SIZE 53.200 BY 765.000 ;
END MAS1929

MACRO MAS1930
     SIZE 29.200 BY 36.000 ;
END MAS1930

MACRO MAS1931
     SIZE 31.500 BY 240.300 ;
END MAS1931

MACRO MAS1933
     SIZE 37.800 BY 225.900 ;
END MAS1933

MACRO MAS1939
     SIZE 7.300 BY 7.200 ;
END MAS1939

MACRO MAS1940
     SIZE 7.300 BY 7.200 ;
END MAS1940

END LIBRARY
