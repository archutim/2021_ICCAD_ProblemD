MACRO MAS5165
     SIZE 295.300 BY 180.000 ;
END MAS5165

MACRO MAS5166
     SIZE 64.400 BY 66.600 ;
END MAS5166

MACRO MAS5167
     SIZE 33.600 BY 33.300 ;
END MAS5167

MACRO MAS5171
     SIZE 133.800 BY 174.600 ;
END MAS5171

MACRO MAS5172
     SIZE 54.600 BY 67.500 ;
END MAS5172

MACRO MAS5173
     SIZE 34.100 BY 36.900 ;
END MAS5173

MACRO MAS5174
     SIZE 245.600 BY 440.100 ;
END MAS5174

MACRO MAS5175
     SIZE 41.600 BY 44.100 ;
END MAS5175

MACRO MAS5176
     SIZE 245.600 BY 440.100 ;
END MAS5176

MACRO MAS5177
     SIZE 557.200 BY 377.100 ;
END MAS5177

MACRO MAS5178
     SIZE 64.600 BY 266.400 ;
END MAS5178

MACRO MAS5179
     SIZE 245.600 BY 440.100 ;
END MAS5179

MACRO MAS5180
     SIZE 54.600 BY 67.500 ;
END MAS5180

MACRO MAS5181
     SIZE 41.600 BY 44.100 ;
END MAS5181

MACRO MAS5182
     SIZE 245.600 BY 440.100 ;
END MAS5182

MACRO MAS5183
     SIZE 54.600 BY 67.500 ;
END MAS5183

MACRO MAS5184
     SIZE 41.600 BY 44.100 ;
END MAS5184

MACRO MAS5185
     SIZE 557.200 BY 377.100 ;
END MAS5185

MACRO MAS5186
     SIZE 64.600 BY 266.400 ;
END MAS5186

MACRO MAS5187
     SIZE 245.600 BY 440.100 ;
END MAS5187

MACRO MAS5188
     SIZE 41.600 BY 44.100 ;
END MAS5188

MACRO MAS5189
     SIZE 245.600 BY 440.100 ;
END MAS5189

MACRO MAS5190
     SIZE 41.600 BY 44.100 ;
END MAS5190

MACRO MAS5191
     SIZE 557.200 BY 377.100 ;
END MAS5191

MACRO MAS5192
     SIZE 64.600 BY 266.400 ;
END MAS5192

MACRO MAS5193
     SIZE 245.600 BY 440.100 ;
END MAS5193

MACRO MAS5194
     SIZE 54.600 BY 67.500 ;
END MAS5194

MACRO MAS5195
     SIZE 41.600 BY 44.100 ;
END MAS5195

MACRO MAS5196
     SIZE 245.600 BY 440.100 ;
END MAS5196

MACRO MAS5197
     SIZE 557.200 BY 377.100 ;
END MAS5197

MACRO MAS5198
     SIZE 64.600 BY 266.400 ;
END MAS5198

MACRO MAS5199
     SIZE 245.600 BY 440.100 ;
END MAS5199

MACRO MAS5200
     SIZE 41.600 BY 44.100 ;
END MAS5200

MACRO MAS5201
     SIZE 245.600 BY 440.100 ;
END MAS5201

MACRO MAS5203
     SIZE 557.200 BY 377.100 ;
END MAS5203

MACRO MAS5204
     SIZE 64.600 BY 266.400 ;
END MAS5204

MACRO MAS5205
     SIZE 41.400 BY 399.600 ;
END MAS5205

MACRO MAS5206
     SIZE 41.600 BY 44.100 ;
END MAS5206

MACRO MAS5207
     SIZE 92.400 BY 431.100 ;
END MAS5207

MACRO MAS5208
     SIZE 23.200 BY 29.700 ;
END MAS5208

MACRO MAS5209
     SIZE 41.400 BY 189.900 ;
END MAS5209

MACRO MAS5210
     SIZE 54.600 BY 67.500 ;
END MAS5210

MACRO MAS5211
     SIZE 34.100 BY 36.900 ;
END MAS5211

MACRO MAS5217
     SIZE 44.100 BY 207.000 ;
END MAS5217

MACRO MAS5220
     SIZE 44.100 BY 207.000 ;
END MAS5220

MACRO MAS5223
     SIZE 574.500 BY 252.000 ;
END MAS5223

MACRO MAS5224
     SIZE 64.400 BY 66.600 ;
END MAS5224

MACRO MAS5225
     SIZE 42.300 BY 40.500 ;
END MAS5225

MACRO MAS5226
     SIZE 574.500 BY 252.000 ;
END MAS5226

MACRO MAS5227
     SIZE 574.500 BY 252.000 ;
END MAS5227

MACRO MAS5228
     SIZE 42.300 BY 40.500 ;
END MAS5228

MACRO MAS5230
     SIZE 574.500 BY 252.000 ;
END MAS5230

MACRO MAS5231
     SIZE 133.800 BY 618.300 ;
END MAS5231

MACRO MAS5232
     SIZE 54.600 BY 68.400 ;
END MAS5232

MACRO MAS5233
     SIZE 41.600 BY 44.100 ;
END MAS5233

MACRO MAS5234
     SIZE 574.500 BY 252.000 ;
END MAS5234

MACRO MAS5235
     SIZE 64.400 BY 66.600 ;
END MAS5235

MACRO MAS5236
     SIZE 42.300 BY 40.500 ;
END MAS5236

MACRO MAS5238
     SIZE 574.500 BY 252.000 ;
END MAS5238

MACRO MAS5239
     SIZE 574.500 BY 252.000 ;
END MAS5239

MACRO MAS5240
     SIZE 64.400 BY 66.600 ;
END MAS5240

MACRO MAS5241
     SIZE 42.300 BY 40.500 ;
END MAS5241

MACRO MAS5242
     SIZE 574.500 BY 252.000 ;
END MAS5242

MACRO MAS5243
     SIZE 42.300 BY 40.500 ;
END MAS5243

MACRO MAS5244
     SIZE 133.800 BY 618.300 ;
END MAS5244

MACRO MAS5245
     SIZE 41.600 BY 44.100 ;
END MAS5245

MACRO MAS5246
     SIZE 22.200 BY 231.300 ;
END MAS5246

MACRO MAS5247
     SIZE 22.200 BY 231.300 ;
END MAS5247

MACRO MAS5252
     SIZE 53.500 BY 198.000 ;
END MAS5252

MACRO MAS5253
     SIZE 54.600 BY 67.500 ;
END MAS5253

MACRO MAS5254
     SIZE 21.700 BY 20.700 ;
END MAS5254

MACRO MAS5255
     SIZE 53.500 BY 198.000 ;
END MAS5255

MACRO MAS5256
     SIZE 54.600 BY 67.500 ;
END MAS5256

MACRO MAS5257
     SIZE 21.700 BY 20.700 ;
END MAS5257

MACRO MAS5258
     SIZE 53.500 BY 198.000 ;
END MAS5258

MACRO MAS5259
     SIZE 21.700 BY 20.700 ;
END MAS5259

MACRO MAS5260
     SIZE 53.500 BY 198.000 ;
END MAS5260

MACRO MAS5261
     SIZE 53.500 BY 198.000 ;
END MAS5261

MACRO MAS5262
     SIZE 34.800 BY 210.600 ;
END MAS5262

MACRO MAS5263
     SIZE 46.000 BY 397.800 ;
END MAS5263

MACRO MAS5264
     SIZE 71.600 BY 81.000 ;
END MAS5264

MACRO MAS5265
     SIZE 23.200 BY 29.700 ;
END MAS5265

MACRO MAS5266
     SIZE 34.800 BY 231.300 ;
END MAS5266

MACRO MAS5290
     SIZE 7.300 BY 7.200 ;
END MAS5290

MACRO MAS5310
     SIZE 7.300 BY 7.200 ;
END MAS5310

END LIBRARY
